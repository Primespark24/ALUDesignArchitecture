-------------------------------------------------
-- Module Name: alu - group designed 
-------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.NUMERIC_STD.all;   

entity alu is
    generic ( N : integer := 32 );
    port (  -- the alu connections to external circuitry:
      -- TODO - Design your groups ALU inputs and outputs!
    );-- operation result
end alu;

architecture behavioral of alu is


-- TODO - Design your group's ALU



end behavioral;